fft_pll_inst : fft_pll PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
